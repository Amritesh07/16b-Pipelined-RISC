library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.all;
use work.components.all;

entity Datapath is
end Datapath;

architecture arch of Datapath is

begin




end arch;